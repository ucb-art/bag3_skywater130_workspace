.INCLUDE /mnt/tools/PDK/skywater130_closed/V1.3.0/LVS/Calibre/source.cdl

*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM



.SUBCKT nmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nlowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B plowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phighvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS


.SUBCKT skywater_diffamp v_inn v_inp v_out VDD VSS
*.PININFO v_inn:I v_inp:I v_out:O VDD:B VSS:B
XGMn_left VSS tail_g v_inp tail_n / nmos4_standard l=150n nf=2 w=420n
XGMn_right VSS v_out v_inn tail_n / nmos4_standard l=150n nf=2 w=420n
XGMp_left VDD tail_g v_inp tail_p / pmos4_standard l=150n nf=12 w=550n
XGMp_right VDD v_out v_inn tail_p / pmos4_standard l=150n nf=12 w=550n
XTailn VSS tail_n tail_g VSS / nmos4_standard l=150n nf=4 w=420n
XTailp VDD tail_p tail_g VDD / pmos4_standard l=150n nf=24 w=550n
.ENDS
