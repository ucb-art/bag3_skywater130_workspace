.INCLUDE /mnt/tools/PDK/skywater130_closed/V1.3.0/LVS/Calibre/source.cdl

*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM



.SUBCKT nmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nhvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nlowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT nmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B nshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hv B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phv l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvesd B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phvesd l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_svt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_lvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B plowvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_hvt B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B phighvt l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS

.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
MM0 D G S B pshort l=l*1.0e6 w=w*1.0e6 m=nf mult=1
.ENDS


.SUBCKT skywater_nor2_pmos4_standard_stack2_w110_l30_seg2 b d g<1> g<0> s
*.PININFO b:B d:B g<1>:B g<0>:B s:B
XP_1 b m<1> g<0> s / pmos4_standard l=150n nf=1 w=550n
XP_0 b m<0> g<0> s / pmos4_standard l=150n nf=1 w=550n
XP_3 b d g<1> m<1> / pmos4_standard l=150n nf=1 w=550n
XP_2 b d g<1> m<0> / pmos4_standard l=150n nf=1 w=550n
.ENDS


.SUBCKT skywater_nor2_nmos4_standard_w84_l30_seg1 b d g s
*.PININFO b:B d:B g:B s:B
XN b d g s / nmos4_standard l=150n nf=1 w=420n
.ENDS


.SUBCKT skywater_nor2 in<1> in<0> out VDD VSS
*.PININFO in<1>:I in<0>:I out:O VDD:B VSS:B
XN_1 VSS out in<1> VSS / skywater_nor2_nmos4_standard_w84_l30_seg1
XN_0 VSS out in<0> VSS / skywater_nor2_nmos4_standard_w84_l30_seg1
XP VDD out in<1> in<0> VDD / skywater_nor2_pmos4_standard_stack2_w110_l30_seg2
.ENDS
